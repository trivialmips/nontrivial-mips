`include "cpu_defs.svh"

module cpu_core(
	input  logic       clk,
	input  logic       rst_n,
	cpu_ibus_if.master ibus,
	cpu_dbus_if.master dbus
);

endmodule
