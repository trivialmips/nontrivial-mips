`ifndef CPU_DEFS_SVH
`define CPU_DEFS_SVH

/*
	This header defines data structures and constants used in CPU internally
*/

`endif
