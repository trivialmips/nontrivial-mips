// this file is only a Verilog wrapper of NonTrivialMIPS CPU in SoC block design
// for SystemVerilog file cannot be used as modules in BDs

module nontrivial_mips #(
	parameter BUS_WIDTH = 4
) (
    // external signals
    input  wire        aclk   ,
    input  wire        reset_n,
    input  wire [4 :0] intr   ,

    // icache
	// AXI AR signals
	output wire [BUS_WIDTH - 1 :0] icache_arid   ,
	output wire [31:0]             icache_araddr ,
	output wire [3 :0]             icache_arlen  ,
	output wire [2 :0]             icache_arsize ,
	output wire [1 :0]             icache_arburst,
	output wire [1 :0]             icache_arlock ,
	output wire [3 :0]             icache_arcache,
	output wire [2 :0]             icache_arprot ,
	output wire                    icache_arvalid,
	input  wire                    icache_arready,
	// AXI R signals
	input  wire [BUS_WIDTH - 1 :0] icache_rid    ,
	input  wire [31:0]             icache_rdata  ,
	input  wire [1 :0]             icache_rresp  ,
	input  wire                    icache_rlast  ,
	input  wire                    icache_rvalid ,
	output wire                    icache_rready ,
	// AXI AW signals
	output wire [BUS_WIDTH - 1 :0] icache_awid   ,
	output wire [31:0]             icache_awaddr ,
	output wire [3 :0]             icache_awlen  ,
	output wire [2 :0]             icache_awsize ,
	output wire [1 :0]             icache_awburst,
	output wire [1 :0]             icache_awlock ,
	output wire [3 :0]             icache_awcache,
	output wire [2 :0]             icache_awprot ,
	output wire                    icache_awvalid,
	input  wire                    icache_awready,
	// AXI W signals
	output wire [BUS_WIDTH - 1 :0] icache_wid    ,
	output wire [31:0]             icache_wdata  ,
	output wire [3 :0]             icache_wstrb  ,
	output wire                    icache_wlast  ,
	output wire                    icache_wvalid ,
	input  wire                    icache_wready ,
	// AXI B signals
	input  wire [BUS_WIDTH - 1 :0] icache_bid    ,
	input  wire [1 :0]             icache_bresp  ,
	input  wire                    icache_bvalid ,
	output wire                    icache_bready ,

    // dcache
	// AXI AR signals
	output wire [BUS_WIDTH - 1 :0] dcache_arid   ,
	output wire [31:0]             dcache_araddr ,
	output wire [3 :0]             dcache_arlen  ,
	output wire [2 :0]             dcache_arsize ,
	output wire [1 :0]             dcache_arburst,
	output wire [1 :0]             dcache_arlock ,
	output wire [3 :0]             dcache_arcache,
	output wire [2 :0]             dcache_arprot ,
	output wire                    dcache_arvalid,
	input  wire                    dcache_arready,
	// AXI R signals
	input  wire [BUS_WIDTH - 1 :0] dcache_rid    ,
	input  wire [31:0]             dcache_rdata  ,
	input  wire [1 :0]             dcache_rresp  ,
	input  wire                    dcache_rlast  ,
	input  wire                    dcache_rvalid ,
	output wire                    dcache_rready ,
	// AXI AW signals
	output wire [BUS_WIDTH - 1 :0] dcache_awid   ,
	output wire [31:0]             dcache_awaddr ,
	output wire [3 :0]             dcache_awlen  ,
	output wire [2 :0]             dcache_awsize ,
	output wire [1 :0]             dcache_awburst,
	output wire [1 :0]             dcache_awlock ,
	output wire [3 :0]             dcache_awcache,
	output wire [2 :0]             dcache_awprot ,
	output wire                    dcache_awvalid,
	input  wire                    dcache_awready,
	// AXI W signals
	output wire [BUS_WIDTH - 1 :0] dcache_wid    ,
	output wire [31:0]             dcache_wdata  ,
	output wire [3 :0]             dcache_wstrb  ,
	output wire                    dcache_wlast  ,
	output wire                    dcache_wvalid ,
	input  wire                    dcache_wready ,
	// AXI B signals
	input  wire [BUS_WIDTH - 1 :0] dcache_bid    ,
	input  wire [1 :0]             dcache_bresp  ,
	input  wire                    dcache_bvalid ,
	output wire                    dcache_bready ,

	// uncached
	// AXI AR signals
	output wire [BUS_WIDTH - 1 :0] uncached_arid   ,
	output wire [31:0]             uncached_araddr ,
	output wire [3 :0]             uncached_arlen  ,
	output wire [2 :0]             uncached_arsize ,
	output wire [1 :0]             uncached_arburst,
	output wire [1 :0]             uncached_arlock ,
	output wire [3 :0]             uncached_arcache,
	output wire [2 :0]             uncached_arprot ,
	output wire                    uncached_arvalid,
	input  wire                    uncached_arready,
	// AXI R signals
	input  wire [BUS_WIDTH - 1 :0] uncached_rid    ,
	input  wire [31:0]             uncached_rdata  ,
	input  wire [1 :0]             uncached_rresp  ,
	input  wire                    uncached_rlast  ,
	input  wire                    uncached_rvalid ,
	output wire                    uncached_rready ,
	// AXI AW signals
	output wire [BUS_WIDTH - 1 :0] uncached_awid   ,
	output wire [31:0]             uncached_awaddr ,
	output wire [3 :0]             uncached_awlen  ,
	output wire [2 :0]             uncached_awsize ,
	output wire [1 :0]             uncached_awburst,
	output wire [1 :0]             uncached_awlock ,
	output wire [3 :0]             uncached_awcache,
	output wire [2 :0]             uncached_awprot ,
	output wire                    uncached_awvalid,
	input  wire                    uncached_awready,
	// AXI W signals
	output wire [BUS_WIDTH - 1 :0] uncached_wid    ,
	output wire [31:0]             uncached_wdata  ,
	output wire [3 :0]             uncached_wstrb  ,
	output wire                    uncached_wlast  ,
	output wire                    uncahced_wvalid ,
	input  wire                    uncached_wready ,
	// AXI B signals
	input  wire [BUS_WIDTH - 1 :0] uncached_bid    ,
	input  wire [1 :0]             uncached_bresp  ,
	input  wire                    uncached_bvalid ,
	output wire                    uncached_bready
);

    // connect all signals as-is
    nontrivial_mips_impl cpu_impl(
        .aclk            (aclk            ),
        .reset_n         (reset_n         ),
        .intr            (intr            ),
        .icache_arid     (icache_arid     ),
        .icache_araddr   (icache_araddr   ),
        .icache_arlen    (icache_arlen    ),
        .icache_arsize   (icache_arsize   ),
        .icache_arburst  (icache_arburst  ),
        .icache_arlock   (icache_arlock   ),
        .icache_arcache  (icache_arcache  ),
        .icache_arprot   (icache_arprot   ),
        .icache_arvalid  (icache_arvalid  ),
        .icache_arready  (icache_arready  ),
        .icache_rid      (icache_rid      ),
        .icache_rdata    (icache_rdata    ),
        .icache_rresp    (icache_rresp    ),
        .icache_rlast    (icache_rlast    ),
        .icache_rvalid   (icache_rvalid   ),
        .icache_rready   (icache_rready   ),
        .icache_awid     (icache_awid     ),
        .icache_awaddr   (icache_awaddr   ),
        .icache_awlen    (icache_awlen    ),
        .icache_awsize   (icache_awsize   ),
        .icache_awburst  (icache_awburst  ),
        .icache_awlock   (icache_awlock   ),
        .icache_awcache  (icache_awcache  ),
        .icache_awprot   (icache_awprot   ),
        .icache_awvalid  (icache_awvalid  ),
        .icache_awready  (icache_awready  ),
        .icache_wid      (icache_wid      ),
        .icache_wdata    (icache_wdata    ),
        .icache_wstrb    (icache_wstrb    ),
        .icache_wlast    (icache_wlast    ),
        .icache_wvalid   (icache_wvalid   ),
        .icache_wready   (icache_wready   ),
        .icache_bid      (icache_bid      ),
        .icache_bresp    (icache_bresp    ),
        .icache_bvalid   (icache_bvalid   ),
        .icache_bready   (icache_bready   ),
        .dcache_arid     (dcache_arid     ),
        .dcache_araddr   (dcache_araddr   ),
        .dcache_arlen    (dcache_arlen    ),
        .dcache_arsize   (dcache_arsize   ),
        .dcache_arburst  (dcache_arburst  ),
        .dcache_arlock   (dcache_arlock   ),
        .dcache_arcache  (dcache_arcache  ),
        .dcache_arprot   (dcache_arprot   ),
        .dcache_arvalid  (dcache_arvalid  ),
        .dcache_arready  (dcache_arready  ),
        .dcache_rid      (dcache_rid      ),
        .dcache_rdata    (dcache_rdata    ),
        .dcache_rresp    (dcache_rresp    ),
        .dcache_rlast    (dcache_rlast    ),
        .dcache_rvalid   (dcache_rvalid   ),
        .dcache_rready   (dcache_rready   ),
        .dcache_awid     (dcache_awid     ),
        .dcache_awaddr   (dcache_awaddr   ),
        .dcache_awlen    (dcache_awlen    ),
        .dcache_awsize   (dcache_awsize   ),
        .dcache_awburst  (dcache_awburst  ),
        .dcache_awlock   (dcache_awlock   ),
        .dcache_awcache  (dcache_awcache  ),
        .dcache_awprot   (dcache_awprot   ),
        .dcache_awvalid  (dcache_awvalid  ),
        .dcache_awready  (dcache_awready  ),
        .dcache_wid      (dcache_wid      ),
        .dcache_wdata    (dcache_wdata    ),
        .dcache_wstrb    (dcache_wstrb    ),
        .dcache_wlast    (dcache_wlast    ),
        .dcache_wvalid   (dcache_wvalid   ),
        .dcache_wready   (dcache_wready   ),
        .dcache_bid      (dcache_bid      ),
        .dcache_bresp    (dcache_bresp    ),
        .dcache_bvalid   (dcache_bvalid   ),
        .dcache_bready   (dcache_bready   ),
        .uncached_arid   (uncached_arid   ),
        .uncached_araddr (uncached_araddr ),
        .uncached_arlen  (uncached_arlen  ),
        .uncached_arsize (uncached_arsize ),
        .uncached_arburst(uncached_arburst),
        .uncached_arlock (uncached_arlock ),
        .uncached_arcache(uncached_arcache),
        .uncached_arprot (uncached_arprot ),
        .uncached_arvalid(uncached_arvalid),
        .uncached_arready(uncached_arready),
        .uncached_rid    (uncached_rid    ),
        .uncached_rdata  (uncached_rdata  ),
        .uncached_rresp  (uncached_rresp  ),
        .uncached_rlast  (uncached_rlast  ),
        .uncached_rvalid (uncached_rvalid ),
        .uncached_rready (uncached_rready ),
        .uncached_awid   (uncached_awid   ),
        .uncached_awaddr (uncached_awaddr ),
        .uncached_awlen  (uncached_awlen  ),
        .uncached_awsize (uncached_awsize ),
        .uncached_awburst(uncached_awburst),
        .uncached_awlock (uncached_awlock ),
        .uncached_awcache(uncached_awcache),
        .uncached_awprot (uncached_awprot ),
        .uncached_awvalid(uncached_awvalid),
        .uncached_awready(uncached_awready),
        .uncached_wid    (uncached_wid    ),
        .uncached_wdata  (uncached_wdata  ),
        .uncached_wstrb  (uncached_wstrb  ),
        .uncached_wlast  (uncached_wlast  ),
        .uncahced_wvalid (uncahced_wvalid ),
        .uncached_wready (uncached_wready ),
        .uncached_bid    (uncached_bid    ),
        .uncached_bresp  (uncached_bresp  ),
        .uncached_bvalid (uncached_bvalid ),
        .uncached_bready (uncached_bready )
    );

endmodule
