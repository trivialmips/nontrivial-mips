`ifndef CACHE_DEFS_SVH
`define CACHE_DEFS_SVH

`endif
