`include "cpu_defs.svh"

module instr_queue(
	input  logic clk,
	input  logic rst_n
);

endmodule
