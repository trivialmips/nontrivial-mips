`ifndef COMPILE_OPTIONS_SVH
`define COMPILE_OPTIONS_SVH

/**
    Options to control optional components to be compiled
    These options are used to speed up compilation when debugging

**/

`define CPU_MMU_ENABLED 1
`define CPU_CP0_ENABLED 1
`define CPU_CP1_ENABLED 1
`define CPU_SUPERSCALAR_ENABLED 1

`endif
