`include "cpu_defs.svh"

module nontrivial_mips(
	input  logic       clk,
	input  logic       rst_n,
	cpu_ibus_if.master ibus,
	cpu_dbus_if.master dbus
);

endmodule
