// this file is only a Verilog wrapper of NonTrivialMIPS CPU
// for SystemVerilog file cannot be used as modules in block design

module nontrivial_mips #(
	parameter BUS_WIDTH = 4
) (
    // external signals
    input  wire [4 :0] intr   ,
    input  wire        aclk   ,
    input  wire        reset_n,

    // icache
	// AXI AR signals
	output wire [BUS_WIDTH - 1 :0] arid_icache   ,
	output wire [31:0]             araddr_icache ,
	output wire [3 :0]             arlen_icache  ,
	output wire [2 :0]             arsize_icache ,
	output wire [1 :0]             arburst_icache,
	output wire [1 :0]             arlock_icache ,
	output wire [3 :0]             arcache_icache,
	output wire [2 :0]             arprot_icache ,
	output wire                    arvalid_icache,
	input  wire                    arready_icache,
	// AXI R signals
	input  wire [BUS_WIDTH - 1 :0] rid_icache    ,
	input  wire [31:0]             rdata_icache  ,
	input  wire [1 :0]             rresp_icache  ,
	input  wire                    rlast_icache  ,
	input  wire                    rvalid_icache ,
	output wire                    rready_icache ,
	// AXI AW signals
	output wire [BUS_WIDTH - 1 :0] awid_icache   ,
	output wire [31:0]             awaddr_icache ,
	output wire [3 :0]             awlen_icache  ,
	output wire [2 :0]             awsize_icache ,
	output wire [1 :0]             awburst_icache,
	output wire [1 :0]             awlock_icache ,
	output wire [3 :0]             awcache_icache,
	output wire [2 :0]             awprot_icache ,
	output wire                    awvalid_icache,
	input  wire                    awready_icache,
	// AXI W signals
	output wire [BUS_WIDTH - 1 :0] wid_icache    ,
	output wire [31:0]             wdata_icache  ,
	output wire [3 :0]             wstrb_icache  ,
	output wire                    wlast_icache  ,
	output wire                    wvalid_icache ,
	input  wire                    wready_icache ,
	// AXI B signals
	input  wire [BUS_WIDTH - 1 :0] bid_icache    ,
	input  wire [1 :0]             bresp_icache  ,
	input  wire                    bvalid_icache ,
	output wire                    bready_icache ,

    // dcache
	// AXI AR signals
	output wire [BUS_WIDTH - 1 :0] arid_dcache   ,
	output wire [31:0]             araddr_dcache ,
	output wire [3 :0]             arlen_dcache  ,
	output wire [2 :0]             arsize_dcache ,
	output wire [1 :0]             arburst_dcache,
	output wire [1 :0]             arlock_dcache ,
	output wire [3 :0]             arcache_dcache,
	output wire [2 :0]             arprot_dcache ,
	output wire                    arvalid_dcache,
	input  wire                    arready_dcache,
	// AXI R signals
	input  wire [BUS_WIDTH - 1 :0] rid_dcache    ,
	input  wire [31:0]             rdata_dcache  ,
	input  wire [1 :0]             rresp_dcache  ,
	input  wire                    rlast_dcache  ,
	input  wire                    rvalid_dcache ,
	output wire                    rready_dcache ,
	// AXI AW signals
	output wire [BUS_WIDTH - 1 :0] awid_dcache   ,
	output wire [31:0]             awaddr_dcache ,
	output wire [3 :0]             awlen_dcache  ,
	output wire [2 :0]             awsize_dcache ,
	output wire [1 :0]             awburst_dcache,
	output wire [1 :0]             awlock_dcache ,
	output wire [3 :0]             awcache_dcache,
	output wire [2 :0]             awprot_dcache ,
	output wire                    awvalid_dcache,
	input  wire                    awready_dcache,
	// AXI W signals
	output wire [BUS_WIDTH - 1 :0] wid_dcache    ,
	output wire [31:0]             wdata_dcache  ,
	output wire [3 :0]             wstrb_dcache  ,
	output wire                    wlast_dcache  ,
	output wire                    wvalid_dcache ,
	input  wire                    wready_dcache ,
	// AXI B signals
	input  wire [BUS_WIDTH - 1 :0] bid_dcache    ,
	input  wire [1 :0]             bresp_dcache  ,
	input  wire                    bvalid_dcache ,
	output wire                    bready_dcache
);

    // negate the polarity of reset signal
    wire reset = ~reset_n;

    // connect all signals as-is
    nontrivial_mips_impl cpu_impl(
        .intr          (intr          ),
        .aclk          (aclk          ),
        .reset_n       (reset_n       ),
        .arid_icache   (arid_icache   ),
        .araddr_icache (araddr_icache ),
        .arlen_icache  (arlen_icache  ),
        .arsize_icache (arsize_icache ),
        .arburst_icache(arburst_icache),
        .arlock_icache (arlock_icache ),
        .arcache_icache(arcache_icache),
        .arprot_icache (arprot_icache ),
        .arvalid_icache(arvalid_icache),
        .arready_icache(arready_icache),
        .rid_icache    (rid_icache    ),
        .rdata_icache  (rdata_icache  ),
        .rresp_icache  (rresp_icache  ),
        .rlast_icache  (rlast_icache  ),
        .rvalid_icache (rvalid_icache ),
        .rready_icache (rready_icache ),
        .awid_icache   (awid_icache   ),
        .awaddr_icache (awaddr_icache ),
        .awlen_icache  (awlen_icache  ),
        .awsize_icache (awsize_icache ),
        .awburst_icache(awburst_icache),
        .awlock_icache (awlock_icache ),
        .awcache_icache(awcache_icache),
        .awprot_icache (awprot_icache ),
        .awvalid_icache(awvalid_icache),
        .awready_icache(awready_icache),
        .wid_icache    (wid_icache    ),
        .wdata_icache  (wdata_icache  ),
        .wstrb_icache  (wstrb_icache  ),
        .wlast_icache  (wlast_icache  ),
        .wvalid_icache (wvalid_icache ),
        .wready_icache (wready_icache ),
        .bid_icache    (bid_icache    ),
        .bresp_icache  (bresp_icache  ),
        .bvalid_icache (bvalid_icache ),
        .bready_icache (bready_icache ),
        .arid_dcache   (arid_dcache   ),
        .araddr_dcache (araddr_dcache ),
        .arlen_dcache  (arlen_dcache  ),
        .arsize_dcache (arsize_dcache ),
        .arburst_dcache(arburst_dcache),
        .arlock_dcache (arlock_dcache ),
        .arcache_dcache(arcache_dcache),
        .arprot_dcache (arprot_dcache ),
        .arvalid_dcache(arvalid_dcache),
        .arready_dcache(arready_dcache),
        .rid_dcache    (rid_dcache    ),
        .rdata_dcache  (rdata_dcache  ),
        .rresp_dcache  (rresp_dcache  ),
        .rlast_dcache  (rlast_dcache  ),
        .rvalid_dcache (rvalid_dcache ),
        .rready_dcache (rready_dcache ),
        .awid_dcache   (awid_dcache   ),
        .awaddr_dcache (awaddr_dcache ),
        .awlen_dcache  (awlen_dcache  ),
        .awsize_dcache (awsize_dcache ),
        .awburst_dcache(awburst_dcache),
        .awlock_dcache (awlock_dcache ),
        .awcache_dcache(awcache_dcache),
        .awprot_dcache (awprot_dcache ),
        .awvalid_dcache(awvalid_dcache),
        .awready_dcache(awready_dcache),
        .wid_dcache    (wid_dcache    ),
        .wdata_dcache  (wdata_dcache  ),
        .wstrb_dcache  (wstrb_dcache  ),
        .wlast_dcache  (wlast_dcache  ),
        .wvalid_dcache (wvalid_dcache ),
        .wready_dcache (wready_dcache ),
        .bid_dcache    (bid_dcache    ),
        .bresp_dcache  (bresp_dcache  ),
        .bvalid_dcache (bvalid_dcache ),
        .bready_dcache (bready_dcache )
    );

endmodule
