`include "cpu_defs.svh"

module alu(
);

endmodule
