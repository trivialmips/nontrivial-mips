`include "cpu_defs.svh"

module instr_exec #(
	parameter int ALU_SIZE = 4
) (
	input  logic         clk,
	input  logic         rst
);

endmodule
