`ifndef COMPILE_OPTION_SVH
`define COMPILE_OPTION_SVH

/*
    Options to control optional components to be compiled
    These options are used to speed up compilation when debugging

*/


`endif
